module mux_5_x_32_decoder (select, out);
parameter n = 64;
parameter log_2_n = log2(n);
input  [log_2_n-1:0] select;
output [n-1:0] out;

reg [n-1:0] out_reg;

always begin
    case(select)
        5'd00 : out_reg <= 64'b00000000000000000000000000000001;
        5'd01 : out_reg <= 64'b00000000000000000000000000000010;
        5'd02 : out_reg <= 64'b00000000000000000000000000000100;
        5'd03 : out_reg <= 64'b00000000000000000000000000001000;
        5'd04 : out_reg <= 64'b00000000000000000000000000010000;
        5'd05 : out_reg <= 64'b00000000000000000000000000100000;
        5'd06 : out_reg <= 64'b00000000000000000000000001000000;
        5'd07 : out_reg <= 64'b00000000000000000000000010000000;
        5'd08 : out_reg <= 64'b00000000000000000000000100000000;
        5'd09 : out_reg <= 64'b00000000000000000000001000000000;
        5'd10 : out_reg <= 64'b00000000000000000000010000000000;
        5'd11 : out_reg <= 64'b00000000000000000000100000000000;
        5'd12 : out_reg <= 64'b00000000000000000001000000000000;
        5'd13 : out_reg <= 64'b00000000000000000010000000000000;
        5'd14 : out_reg <= 64'b00000000000000000100000000000000;
        5'd15 : out_reg <= 64'b00000000000000001000000000000000;
        5'd16 : out_reg <= 64'b00000000000000010000000000000000;
        5'd17 : out_reg <= 64'b00000000000000100000000000000000;
        5'd18 : out_reg <= 64'b00000000000001000000000000000000;
        5'd19 : out_reg <= 64'b00000000000010000000000000000000;
        5'd20 : out_reg <= 64'b00000000000100000000000000000000;
        5'd21 : out_reg <= 64'b00000000001000000000000000000000;
        5'd22 : out_reg <= 64'b00000000010000000000000000000000;
        5'd23 : out_reg <= 64'b00000000100000000000000000000000;
        5'd24 : out_reg <= 64'b00000001000000000000000000000000;
        5'd25 : out_reg <= 64'b00000010000000000000000000000000;
        5'd26 : out_reg <= 64'b00000100000000000000000000000000;
        5'd27 : out_reg <= 64'b00001000000000000000000000000000;
        5'd28 : out_reg <= 64'b00010000000000000000000000000000;
        5'd29 : out_reg <= 64'b00100000000000000000000000000000;
        5'd30 : out_reg <= 64'b01000000000000000000000000000000;
        5'd31 : out_reg <= 64'b10000000000000000000000000000000;
    endcase
end

assign out = out_reg;

function log2;
    input x;
    reg i, log;
    begin
        i = x;
        log = 1;
        while(i!=1) begin
            i=i/2;
            log = log + 1;
        end
    end
endfunction

endmodule
