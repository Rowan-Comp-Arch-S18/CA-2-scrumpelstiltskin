module VGA_Testbench();

    reg clk;
    wire [3:0] red_out, green_out, blue_out;
    wire h_sync_out, v_sync_out;

    wire [11:0] h_position;
    wire [10:0] v_position;
    wire [10:0] pixel_position;

    wire out;

    reg [1200:0] data;

    initial begin
        data[39:0]      <= 40'b1010101010101010101010101010101010101010;
        data[79:40]     <= 40'b0101010101010101010101010101010101010101;
        data[119:80]    <= 40'b1010101010101010101010101010101010101010;
        data[159:120]   <= 40'b0101010101010101010101010101010101010101;
        data[199:160]   <= 40'b1010101010101010101010101010101010101010;
        data[239:200]   <= 40'b0101010101010101010101010101010101010101;
        data[279:240]   <= 40'b1010101010101010101010101010101010101010;
        data[319:280]   <= 40'b0101010101010101010101010101010101010101;
        data[359:320]   <= 40'b1010101010101010101010101010101010101010;
        data[399:360]   <= 40'b0101010101010101010101010101010101010101;
        data[439:400]   <= 40'b1010101010101010101010101010101010101010;
        data[479:440]   <= 40'b0101010101010101010101010101010101010101;
        data[519:480]   <= 40'b1010101010101010101010101010101010101010;
        data[559:520]   <= 40'b0101010101010101010101010101010101010101;
        data[599:560]   <= 40'b1010101010101010101010101010101010101010;
        data[639:600]   <= 40'b0101010101010101010101010101010101010101;
        data[679:640]   <= 40'b1010101010101010101010101010101010101010;
        data[719:680]   <= 40'b0101010101010101010101010101010101010101;
        data[759:720]   <= 40'b1010101010101010101010101010101010101010;
        data[799:760]   <= 40'b0101010101010101010101010101010101010101;
        data[839:800]   <= 40'b1010101010101010101010101010101010101010;
        data[879:840]   <= 40'b0101010101010101010101010101010101010101;
        data[919:880]   <= 40'b1010101010101010101010101010101010101010;
        data[959:920]   <= 40'b0101010101010101010101010101010101010101;
        data[999:960]   <= 40'b1010101010101010101010101010101010101010;
        data[1039:1000] <= 40'b0101010101010101010101010101010101010101;
        data[1079:1040] <= 40'b1010101010101010101010101010101010101010;
        data[1119:1080] <= 40'b0101010101010101010101010101010101010101;
        data[1159:1120] <= 40'b1010101010101010101010101010101010101010;
        data[1199:1160] <= 40'b0101010101010101010101010101010101010101;
    end

    VGA_Test vga (
        clk,
        data,
        red_out,
        green_out,
        blue_out,
        h_sync_out,
        v_sync_out,
        h_position,
        v_position,
        pixel_position,
        out
    );

    initial begin
        clk <= 1'b0;
    end

    always begin
        #10000 clk <= ~clk;
    end

    always begin
        #4000000000 $stop;
    end

endmodule

