module mouse_testbench();

			reg PS2_data;
			reg PS2_clk;
			reg system_clk;
			reg reset;
			
			