module program_counter(ps, in, pc);
    // PS
    // 00 PC <- PC
    // 01 PC <- PC + 4
    //
