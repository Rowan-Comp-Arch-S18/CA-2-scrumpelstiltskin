module keyboard(PS2_data, PS2_clk, system_clk, data);

    input PS2_data;
    input PS2_clk;
    input system_clk;

    output [63:0] data;


    registerfile

endmodule
